	end if;
	end process reset_values;

end architecture RTL;

